/*** 
 * @Author: jia200151@126.com
 * @Date: 2025-11-29 10:40:19
 * @LastEditors: lwj
 * @LastEditTime: 2025-11-29 10:44:06
 * @FilePath: \rtl\Neural_engine\conv.v
 * @Description: 
 * @Copyright (c) 2025 by lwj email: jia200151@126.com, All Rights Reserved.
 */
module conv (
    
);
    
endmodule
