/*** 
 * @Author: jia200151@126.com
 * @Date: 2025-12-29 14:51:04
 * @LastEditors: lwj
 * @LastEditTime: 2026-01-09 17:08:05
 * @FilePath: \core\core_controller.v
 * @Description: 
 * @Copyright (c) 2025 by lwj email: jia200151@126.com, All Rights Reserved.
 */
module core_controller (
    input wire clk,
    input wire reset,
    input wire start,
    
    // Control Signals
    input reg decoded_ret,

    // Memory Access State
    input reg [2:0] fetcher_state,
    input reg [2:0] lsu_state ,

    // Current & Next PC
    output reg [7:0] current_pc,
    input reg [7:0] next_pc ,

    // Execution State
    output reg [2:0] core_state,
    output reg done
);
    localparam IDLE = 3'b000, // Waiting to start
        FETCH = 3'b001,       // Fetch instructions from program memory
        DECODE = 3'b010,      // Decode instructions into control signals
        REQUEST = 3'b011,     // Request data from registers or memory
        WAIT = 3'b100,        // Wait for response from memory if necessary
        EXECUTE = 3'b101,     // Execute ALU and PC calculations
        UPDATE = 3'b110,      // Update registers, NZP, and PC
        DONE = 3'b111;        // Done executing this core
    reg any_lsu_waiting = 1'b0;
    always @(posedge clk) begin 
        if (reset) begin
            current_pc <= 0;
            core_state <= IDLE;
            done <= 0;
            any_lsu_waiting = 1'b0;
        end else begin 
            case (core_state)
                IDLE: begin
                    // Here after reset (before kernel is launched, or after previous block has been processed)
                    if (start) begin 
                        // Start by fetching the next instruction for this block based on PC
                        core_state <= FETCH;
                    end
                end
                FETCH: begin 
                    // Move on once fetcher_state = FETCHED
                    if (fetcher_state == 3'b010) begin 
                        core_state <= DECODE;
                    end
                end
                DECODE: begin
                    // Decode is synchronous so we move on after one cycle
                    core_state <= REQUEST;
                end
                REQUEST: begin 
                    // Request is synchronous so we move on after one cycle
                    core_state <= WAIT;
                end
                WAIT: begin
                    // Wait for all LSUs to finish their request before continuing
                    any_lsu_waiting <= 1'b0;

                        // Make sure no lsu_state = REQUESTING or WAITING
                    if (lsu_state == 2'b01 || lsu_state == 2'b10) begin
                        any_lsu_waiting <= 1'b1;
                    end

                    // If no LSU is waiting for a response, move onto the next stage
                    if (!any_lsu_waiting) begin
                        core_state <= EXECUTE;
                    end
                end
                EXECUTE: begin
                    // Execute is synchronous so we move on after one cycle
                    core_state <= UPDATE;
                end
                UPDATE: begin 
                    if (decoded_ret) begin 
                        // If we reach a RET instruction, this block is done executing
                        done <= 1;
                        core_state <= DONE;
                    end else begin 
                        // TODO: Branch divergence. For now assume all next_pc converge
                        current_pc <= next_pc;

                        // Update is synchronous so we move on after one cycle
                        core_state <= FETCH;
                    end
                end
                DONE: begin 
                    // no-op
                end
            endcase
        end
    end
    
endmodule
